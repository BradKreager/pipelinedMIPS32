module dmem (
         input  wire        clk,
         input  wire        we,
         input  wire [5:0]  a,
         input  wire [31:0] d,
         output wire [31:0] q
       );

reg [31:0] ram [0:63];
reg [5:0] addr;

integer n;

initial
  begin
    for (n = 0; n < 64; n = n + 1)
      ram[n] = 32'hFFFFFFFF;
  end

always @ (posedge clk)
  begin
    if (we)
      ram[a] <= d;
  end

always @ (negedge clk)
  begin
    addr <= a;
  end

assign q = ram[addr];

endmodule
